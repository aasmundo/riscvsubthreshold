library IEEE;
use IEEE.STD_LOGIC_1164.all;
library work;
use work.constants.all;


entity instruction_decode is
	port(
	
	);
end instruction_decode;


architecture behave of instruction_decode is

begin
	
end behave;
