../modules/soc_top_tb_no_startup.vhd